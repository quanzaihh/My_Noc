`timescale 1ns / 1ps
/*
    created by: <Xidian University>
    created date: 2024-05-16
*/

module Noc_connector(
    input                           noc_clk,
    input                           rst_n,    
    input   [0:0]                   Noc_0_0_channel0_receive_valid,
    output  [0:0]                   Noc_0_0_channel0_receive_ready,
    input   [`Noc_Data_Width-1:0]   Noc_0_0_channel0_receive_flit,
    output  [0:0]                   Noc_0_0_channel0_receive_VCready,
    input   [0:0]                   Noc_0_0_channel0_receive_is_header,
    input   [0:0]                   Noc_0_0_channel0_receive_is_tail,             
);
                                                                   
                                                                   
endmodule