`timescale 1ps/1ps

module simulation_top