`timescale 1ns / 1ps
/*
    created by: <Xidian University>
    created date: 2024-05-16
*/

module Noc_bridge(
    input                               noc_clk,
    input                               rst_n,    
    input                   
);
                                                                   
                                                                   
endmodule